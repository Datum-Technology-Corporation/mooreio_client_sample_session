`ifndef DATA_WIDTH
`define DATA_WIDTH 8
`endif